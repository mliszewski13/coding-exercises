`include "quadra.svh"

module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = 22'sh34afb1;
        7'b0000001 :  a = 22'sh350b9a;
        7'b0000010 :  a = 22'sh356a3f;
        7'b0000011 :  a = 22'sh35cb8a;
        7'b0000100 :  a = 22'sh362f63;
        7'b0000101 :  a = 22'sh3695af;
        7'b0000110 :  a = 22'sh36fe56;
        7'b0000111 :  a = 22'sh37693d;
        7'b0001000 :  a = 22'sh37d64a;
        7'b0001001 :  a = 22'sh384561;
        7'b0001010 :  a = 22'sh38b667;
        7'b0001011 :  a = 22'sh39293f;
        7'b0001100 :  a = 22'sh399dcd;
        7'b0001101 :  a = 22'sh3a13f3;
        7'b0001110 :  a = 22'sh3a8b95;
        7'b0001111 :  a = 22'sh3b0493;
        7'b0010000 :  a = 22'sh3b7ed0;
        7'b0010001 :  a = 22'sh3bfa2e;
        7'b0010010 :  a = 22'sh3c768d;
        7'b0010011 :  a = 22'sh3cf3ce;
        7'b0010100 :  a = 22'sh3d71d3;
        7'b0010101 :  a = 22'sh3df07a;
        7'b0010110 :  a = 22'sh3e6fa6;
        7'b0010111 :  a = 22'sh3eef36;
        7'b0011000 :  a = 22'sh3f6f0a;
        7'b0011001 :  a = 22'sh3fef02;
        7'b0011010 :  a = 22'sh006eff;
        7'b0011011 :  a = 22'sh00eee0;
        7'b0011100 :  a = 22'sh016e85;
        7'b0011101 :  a = 22'sh01edce;
        7'b0011110 :  a = 22'sh026c9c;
        7'b0011111 :  a = 22'sh02eacf;
        7'b0100000 :  a = 22'sh036847;
        7'b0100001 :  a = 22'sh03e4e5;
        7'b0100010 :  a = 22'sh04608a;
        7'b0100011 :  a = 22'sh04db17;
        7'b0100100 :  a = 22'sh05546d;
        7'b0100101 :  a = 22'sh05cc6e;
        7'b0100110 :  a = 22'sh0642fc;
        7'b0100111 :  a = 22'sh06b7f9;
        7'b0101000 :  a = 22'sh072b48;
        7'b0101001 :  a = 22'sh079ccd;
        7'b0101010 :  a = 22'sh080c6a;
        7'b0101011 :  a = 22'sh087a04;
        7'b0101100 :  a = 22'sh08e580;
        7'b0101101 :  a = 22'sh094ec2;
        7'b0101110 :  a = 22'sh09b5b1;
        7'b0101111 :  a = 22'sh0a1a32;
        7'b0110000 :  a = 22'sh0a7c2d;
        7'b0110001 :  a = 22'sh0adb89;
        7'b0110010 :  a = 22'sh0b382e;
        7'b0110011 :  a = 22'sh0b9206;
        7'b0110100 :  a = 22'sh0be8f8;
        7'b0110101 :  a = 22'sh0c3cf1;
        7'b0110110 :  a = 22'sh0c8dda;
        7'b0110111 :  a = 22'sh0cdba0;
        7'b0111000 :  a = 22'sh0d262f;
        7'b0111001 :  a = 22'sh0d6d75;
        7'b0111010 :  a = 22'sh0db15f;
        7'b0111011 :  a = 22'sh0df1dd;
        7'b0111100 :  a = 22'sh0e2edf;
        7'b0111101 :  a = 22'sh0e6855;
        7'b0111110 :  a = 22'sh0e9e31;
        7'b0111111 :  a = 22'sh0ed065;
        7'b1000000 :  a = 22'sh0efee6;
        7'b1000001 :  a = 22'sh0f29a6;
        7'b1000010 :  a = 22'sh0f509d;
        7'b1000011 :  a = 22'sh0f73bf;
        7'b1000100 :  a = 22'sh0f9305;
        7'b1000101 :  a = 22'sh0fae66;
        7'b1000110 :  a = 22'sh0fc5db;
        7'b1000111 :  a = 22'sh0fd95f;
        7'b1001000 :  a = 22'sh0fe8ed;
        7'b1001001 :  a = 22'sh0ff481;
        7'b1001010 :  a = 22'sh0ffc17;
        7'b1001011 :  a = 22'sh0fffaf;
        7'b1001100 :  a = 22'sh0fff47;
        7'b1001101 :  a = 22'sh0ffadf;
        7'b1001110 :  a = 22'sh0ff278;
        7'b1001111 :  a = 22'sh0fe615;
        7'b1010000 :  a = 22'sh0fd5b8;
        7'b1010001 :  a = 22'sh0fc166;
        7'b1010010 :  a = 22'sh0fa924;
        7'b1010011 :  a = 22'sh0f8cf8;
        7'b1010100 :  a = 22'sh0f6ce8;
        7'b1010101 :  a = 22'sh0f48fe;
        7'b1010110 :  a = 22'sh0f2141;
        7'b1010111 :  a = 22'sh0ef5bc;
        7'b1011000 :  a = 22'sh0ec679;
        7'b1011001 :  a = 22'sh0e9385;
        7'b1011010 :  a = 22'sh0e5ced;
        7'b1011011 :  a = 22'sh0e22bd;
        7'b1011100 :  a = 22'sh0de504;
        7'b1011101 :  a = 22'sh0da3d2;
        7'b1011110 :  a = 22'sh0d5f38;
        7'b1011111 :  a = 22'sh0d1745;
        7'b1100000 :  a = 22'sh0ccc0d;
        7'b1100001 :  a = 22'sh0c7da2;
        7'b1100010 :  a = 22'sh0c2c18;
        7'b1100011 :  a = 22'sh0bd782;
        7'b1100100 :  a = 22'sh0b7ff7;
        7'b1100101 :  a = 22'sh0b258c;
        7'b1100110 :  a = 22'sh0ac858;
        7'b1100111 :  a = 22'sh0a6871;
        7'b1101000 :  a = 22'sh0a05f1;
        7'b1101001 :  a = 22'sh09a0ef;
        7'b1101010 :  a = 22'sh093985;
        7'b1101011 :  a = 22'sh08cfcc;
        7'b1101100 :  a = 22'sh0863e0;
        7'b1101101 :  a = 22'sh07f5db;
        7'b1101110 :  a = 22'sh0785d8;
        7'b1101111 :  a = 22'sh0713f4;
        7'b1110000 :  a = 22'sh06a04b;
        7'b1110001 :  a = 22'sh062afa;
        7'b1110010 :  a = 22'sh05b41e;
        7'b1110011 :  a = 22'sh053bd5;
        7'b1110100 :  a = 22'sh04c23d;
        7'b1110101 :  a = 22'sh044775;
        7'b1110110 :  a = 22'sh03cb9b;
        7'b1110111 :  a = 22'sh034ece;
        7'b1111000 :  a = 22'sh02d12d;
        7'b1111001 :  a = 22'sh0252d8;
        7'b1111010 :  a = 22'sh01d3ee;
        7'b1111011 :  a = 22'sh015490;
        7'b1111100 :  a = 22'sh00d4dc;
        7'b1111101 :  a = 22'sh0054f3;
        7'b1111110 :  a = 22'sh3fd4f5;
        7'b1111111 :  a = 22'sh3f5501;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = 16'sh2d41;
        7'b0000001 :  b = 16'sh2ea6;
        7'b0000010 :  b = 16'sh2ffe;
        7'b0000011 :  b = 16'sh314b;
        7'b0000100 :  b = 16'sh328b;
        7'b0000101 :  b = 16'sh33bf;
        7'b0000110 :  b = 16'sh34e6;
        7'b0000111 :  b = 16'sh35ff;
        7'b0001000 :  b = 16'sh370b;
        7'b0001001 :  b = 16'sh380a;
        7'b0001010 :  b = 16'sh38fa;
        7'b0001011 :  b = 16'sh39dc;
        7'b0001100 :  b = 16'sh3ab0;
        7'b0001101 :  b = 16'sh3b74;
        7'b0001110 :  b = 16'sh3c2a;
        7'b0001111 :  b = 16'sh3cd1;
        7'b0010000 :  b = 16'sh3d69;
        7'b0010001 :  b = 16'sh3df2;
        7'b0010010 :  b = 16'sh3e6b;
        7'b0010011 :  b = 16'sh3ed4;
        7'b0010100 :  b = 16'sh3f2e;
        7'b0010101 :  b = 16'sh3f78;
        7'b0010110 :  b = 16'sh3fb2;
        7'b0010111 :  b = 16'sh3fdc;
        7'b0011000 :  b = 16'sh3ff6;
        7'b0011001 :  b = 16'sh4000;
        7'b0011010 :  b = 16'sh3ffa;
        7'b0011011 :  b = 16'sh3fe4;
        7'b0011100 :  b = 16'sh3fbe;
        7'b0011101 :  b = 16'sh3f89;
        7'b0011110 :  b = 16'sh3f43;
        7'b0011111 :  b = 16'sh3eed;
        7'b0100000 :  b = 16'sh3e88;
        7'b0100001 :  b = 16'sh3e13;
        7'b0100010 :  b = 16'sh3d8f;
        7'b0100011 :  b = 16'sh3cfb;
        7'b0100100 :  b = 16'sh3c58;
        7'b0100101 :  b = 16'sh3ba6;
        7'b0100110 :  b = 16'sh3ae5;
        7'b0100111 :  b = 16'sh3a16;
        7'b0101000 :  b = 16'sh3937;
        7'b0101001 :  b = 16'sh384b;
        7'b0101010 :  b = 16'sh3750;
        7'b0101011 :  b = 16'sh3648;
        7'b0101100 :  b = 16'sh3532;
        7'b0101101 :  b = 16'sh340e;
        7'b0101110 :  b = 16'sh32de;
        7'b0101111 :  b = 16'sh31a1;
        7'b0110000 :  b = 16'sh3058;
        7'b0110001 :  b = 16'sh2f02;
        7'b0110010 :  b = 16'sh2da1;
        7'b0110011 :  b = 16'sh2c34;
        7'b0110100 :  b = 16'sh2abd;
        7'b0110101 :  b = 16'sh293a;
        7'b0110110 :  b = 16'sh27ad;
        7'b0110111 :  b = 16'sh2617;
        7'b0111000 :  b = 16'sh2477;
        7'b0111001 :  b = 16'sh22cd;
        7'b0111010 :  b = 16'sh211b;
        7'b0111011 :  b = 16'sh1f61;
        7'b0111100 :  b = 16'sh1d9f;
        7'b0111101 :  b = 16'sh1bd6;
        7'b0111110 :  b = 16'sh1a05;
        7'b0111111 :  b = 16'sh182e;
        7'b1000000 :  b = 16'sh1651;
        7'b1000001 :  b = 16'sh146f;
        7'b1000010 :  b = 16'sh1287;
        7'b1000011 :  b = 16'sh109b;
        7'b1000100 :  b = 16'sh0eaa;
        7'b1000101 :  b = 16'sh0cb6;
        7'b1000110 :  b = 16'sh0abf;
        7'b1000111 :  b = 16'sh08c5;
        7'b1001000 :  b = 16'sh06c9;
        7'b1001001 :  b = 16'sh04cb;
        7'b1001010 :  b = 16'sh02cc;
        7'b1001011 :  b = 16'sh00cc;
        7'b1001100 :  b = 16'shfecc;
        7'b1001101 :  b = 16'shfccc;
        7'b1001110 :  b = 16'shfacd;
        7'b1001111 :  b = 16'shf8d0;
        7'b1010000 :  b = 16'shf6d4;
        7'b1010001 :  b = 16'shf4db;
        7'b1010010 :  b = 16'shf2e4;
        7'b1010011 :  b = 16'shf0f0;
        7'b1010100 :  b = 16'shef01;
        7'b1010101 :  b = 16'shed15;
        7'b1010110 :  b = 16'sheb2f;
        7'b1010111 :  b = 16'she94d;
        7'b1011000 :  b = 16'she771;
        7'b1011001 :  b = 16'she59c;
        7'b1011010 :  b = 16'she3cd;
        7'b1011011 :  b = 16'she205;
        7'b1011100 :  b = 16'she044;
        7'b1011101 :  b = 16'shde8c;
        7'b1011110 :  b = 16'shdcdb;
        7'b1011111 :  b = 16'shdb34;
        7'b1100000 :  b = 16'shd996;
        7'b1100001 :  b = 16'shd801;
        7'b1100010 :  b = 16'shd676;
        7'b1100011 :  b = 16'shd4f6;
        7'b1100100 :  b = 16'shd381;
        7'b1100101 :  b = 16'shd216;
        7'b1100110 :  b = 16'shd0b7;
        7'b1100111 :  b = 16'shcf64;
        7'b1101000 :  b = 16'shce1d;
        7'b1101001 :  b = 16'shcce3;
        7'b1101010 :  b = 16'shcbb5;
        7'b1101011 :  b = 16'shca95;
        7'b1101100 :  b = 16'shc981;
        7'b1101101 :  b = 16'shc87c;
        7'b1101110 :  b = 16'shc784;
        7'b1101111 :  b = 16'shc69a;
        7'b1110000 :  b = 16'shc5bf;
        7'b1110001 :  b = 16'shc4f2;
        7'b1110010 :  b = 16'shc434;
        7'b1110011 :  b = 16'shc385;
        7'b1110100 :  b = 16'shc2e5;
        7'b1110101 :  b = 16'shc255;
        7'b1110110 :  b = 16'shc1d4;
        7'b1110111 :  b = 16'shc162;
        7'b1111000 :  b = 16'shc100;
        7'b1111001 :  b = 16'shc0ae;
        7'b1111010 :  b = 16'shc06b;
        7'b1111011 :  b = 16'shc039;
        7'b1111100 :  b = 16'shc016;
        7'b1111101 :  b = 16'shc004;
        7'b1111110 :  b = 16'shc001;
        7'b1111111 :  b = 16'shc00e;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = 8'sh5b;
        7'b0000001 :  c = 8'sh58;
        7'b0000010 :  c = 8'sh55;
        7'b0000011 :  c = 8'sh52;
        7'b0000100 :  c = 8'sh4f;
        7'b0000101 :  c = 8'sh4b;
        7'b0000110 :  c = 8'sh48;
        7'b0000111 :  c = 8'sh45;
        7'b0001000 :  c = 8'sh41;
        7'b0001001 :  c = 8'sh3e;
        7'b0001010 :  c = 8'sh3a;
        7'b0001011 :  c = 8'sh37;
        7'b0001100 :  c = 8'sh33;
        7'b0001101 :  c = 8'sh2f;
        7'b0001110 :  c = 8'sh2c;
        7'b0001111 :  c = 8'sh28;
        7'b0010000 :  c = 8'sh24;
        7'b0010001 :  c = 8'sh20;
        7'b0010010 :  c = 8'sh1c;
        7'b0010011 :  c = 8'sh18;
        7'b0010100 :  c = 8'sh14;
        7'b0010101 :  c = 8'sh10;
        7'b0010110 :  c = 8'sh0d;
        7'b0010111 :  c = 8'sh09;
        7'b0011000 :  c = 8'sh05;
        7'b0011001 :  c = 8'sh01;
        7'b0011010 :  c = 8'shfd;
        7'b0011011 :  c = 8'shf9;
        7'b0011100 :  c = 8'shf5;
        7'b0011101 :  c = 8'shf1;
        7'b0011110 :  c = 8'shed;
        7'b0011111 :  c = 8'she9;
        7'b0100000 :  c = 8'she5;
        7'b0100001 :  c = 8'she1;
        7'b0100010 :  c = 8'shdd;
        7'b0100011 :  c = 8'shd9;
        7'b0100100 :  c = 8'shd5;
        7'b0100101 :  c = 8'shd2;
        7'b0100110 :  c = 8'shce;
        7'b0100111 :  c = 8'shca;
        7'b0101000 :  c = 8'shc7;
        7'b0101001 :  c = 8'shc3;
        7'b0101010 :  c = 8'shc0;
        7'b0101011 :  c = 8'shbc;
        7'b0101100 :  c = 8'shb9;
        7'b0101101 :  c = 8'shb6;
        7'b0101110 :  c = 8'shb2;
        7'b0101111 :  c = 8'shaf;
        7'b0110000 :  c = 8'shac;
        7'b0110001 :  c = 8'sha9;
        7'b0110010 :  c = 8'sha6;
        7'b0110011 :  c = 8'sha3;
        7'b0110100 :  c = 8'sha1;
        7'b0110101 :  c = 8'sh9e;
        7'b0110110 :  c = 8'sh9c;
        7'b0110111 :  c = 8'sh99;
        7'b0111000 :  c = 8'sh97;
        7'b0111001 :  c = 8'sh95;
        7'b0111010 :  c = 8'sh92;
        7'b0111011 :  c = 8'sh90;
        7'b0111100 :  c = 8'sh8f;
        7'b0111101 :  c = 8'sh8d;
        7'b0111110 :  c = 8'sh8b;
        7'b0111111 :  c = 8'sh89;
        7'b1000000 :  c = 8'sh88;
        7'b1000001 :  c = 8'sh87;
        7'b1000010 :  c = 8'sh85;
        7'b1000011 :  c = 8'sh84;
        7'b1000100 :  c = 8'sh83;
        7'b1000101 :  c = 8'sh83;
        7'b1000110 :  c = 8'sh82;
        7'b1000111 :  c = 8'sh81;
        7'b1001000 :  c = 8'sh81;
        7'b1001001 :  c = 8'sh80;
        7'b1001010 :  c = 8'sh80;
        7'b1001011 :  c = 8'sh80;
        7'b1001100 :  c = 8'sh80;
        7'b1001101 :  c = 8'sh80;
        7'b1001110 :  c = 8'sh80;
        7'b1001111 :  c = 8'sh81;
        7'b1010000 :  c = 8'sh81;
        7'b1010001 :  c = 8'sh82;
        7'b1010010 :  c = 8'sh83;
        7'b1010011 :  c = 8'sh84;
        7'b1010100 :  c = 8'sh85;
        7'b1010101 :  c = 8'sh86;
        7'b1010110 :  c = 8'sh87;
        7'b1010111 :  c = 8'sh88;
        7'b1011000 :  c = 8'sh8a;
        7'b1011001 :  c = 8'sh8b;
        7'b1011010 :  c = 8'sh8d;
        7'b1011011 :  c = 8'sh8f;
        7'b1011100 :  c = 8'sh91;
        7'b1011101 :  c = 8'sh93;
        7'b1011110 :  c = 8'sh95;
        7'b1011111 :  c = 8'sh97;
        7'b1100000 :  c = 8'sh9a;
        7'b1100001 :  c = 8'sh9c;
        7'b1100010 :  c = 8'sh9f;
        7'b1100011 :  c = 8'sha1;
        7'b1100100 :  c = 8'sha4;
        7'b1100101 :  c = 8'sha7;
        7'b1100110 :  c = 8'shaa;
        7'b1100111 :  c = 8'shad;
        7'b1101000 :  c = 8'shb0;
        7'b1101001 :  c = 8'shb3;
        7'b1101010 :  c = 8'shb6;
        7'b1101011 :  c = 8'shba;
        7'b1101100 :  c = 8'shbd;
        7'b1101101 :  c = 8'shc0;
        7'b1101110 :  c = 8'shc4;
        7'b1101111 :  c = 8'shc7;
        7'b1110000 :  c = 8'shcb;
        7'b1110001 :  c = 8'shcf;
        7'b1110010 :  c = 8'shd2;
        7'b1110011 :  c = 8'shd6;
        7'b1110100 :  c = 8'shda;
        7'b1110101 :  c = 8'shde;
        7'b1110110 :  c = 8'she2;
        7'b1110111 :  c = 8'she6;
        7'b1111000 :  c = 8'she9;
        7'b1111001 :  c = 8'shed;
        7'b1111010 :  c = 8'shf1;
        7'b1111011 :  c = 8'shf5;
        7'b1111100 :  c = 8'shf9;
        7'b1111101 :  c = 8'shfd;
        7'b1111110 :  c = 8'sh01;
        7'b1111111 :  c = 8'sh05;
        default    :  c = 'x;
    endcase

endmodule
