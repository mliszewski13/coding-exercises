`include "quadra.svh"

module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = 32'shf4afb0cd;
        7'b0000001 :  a = 32'shf50b9983;
        7'b0000010 :  a = 32'shf56a3f45;
        7'b0000011 :  a = 32'shf5cb8a69;
        7'b0000100 :  a = 32'shf62f629c;
        7'b0000101 :  a = 32'shf695aeea;
        7'b0000110 :  a = 32'shf6fe55bf;
        7'b0000111 :  a = 32'shf7693cf3;
        7'b0001000 :  a = 32'shf7d649cc;
        7'b0001001 :  a = 32'shf8456108;
        7'b0001010 :  a = 32'shf8b666e2;
        7'b0001011 :  a = 32'shf9293f18;
        7'b0001100 :  a = 32'shf99dccf5;
        7'b0001101 :  a = 32'shfa13f356;
        7'b0001110 :  a = 32'shfa8b94b3;
        7'b0001111 :  a = 32'shfb049323;
        7'b0010000 :  a = 32'shfb7ed068;
        7'b0010001 :  a = 32'shfbfa2df2;
        7'b0010010 :  a = 32'shfc768cec;
        7'b0010011 :  a = 32'shfcf3ce3e;
        7'b0010100 :  a = 32'shfd71d298;
        7'b0010101 :  a = 32'shfdf07a7a;
        7'b0010110 :  a = 32'shfe6fa63b;
        7'b0010111 :  a = 32'shfeef3610;
        7'b0011000 :  a = 32'shff6f0a16;
        7'b0011001 :  a = 32'shffef0259;
        7'b0011010 :  a = 32'sh006efedb;
        7'b0011011 :  a = 32'sh00eedf9e;
        7'b0011100 :  a = 32'sh016e84ab;
        7'b0011101 :  a = 32'sh01edce18;
        7'b0011110 :  a = 32'sh026c9c14;
        7'b0011111 :  a = 32'sh02eaceed;
        7'b0100000 :  a = 32'sh03684715;
        7'b0100001 :  a = 32'sh03e4e531;
        7'b0100010 :  a = 32'sh04608a18;
        7'b0100011 :  a = 32'sh04db16e2;
        7'b0100100 :  a = 32'sh05546cee;
        7'b0100101 :  a = 32'sh05cc6de5;
        7'b0100110 :  a = 32'sh0642fbc8;
        7'b0100111 :  a = 32'sh06b7f8f5;
        7'b0101000 :  a = 32'sh072b482d;
        7'b0101001 :  a = 32'sh079ccc9c;
        7'b0101010 :  a = 32'sh080c69e2;
        7'b0101011 :  a = 32'sh087a0419;
        7'b0101100 :  a = 32'sh08e57fd9;
        7'b0101101 :  a = 32'sh094ec246;
        7'b0101110 :  a = 32'sh09b5b10e;
        7'b0101111 :  a = 32'sh0a1a3277;
        7'b0110000 :  a = 32'sh0a7c2d61;
        7'b0110001 :  a = 32'sh0adb894e;
        7'b0110010 :  a = 32'sh0b382e66;
        7'b0110011 :  a = 32'sh0b920582;
        7'b0110100 :  a = 32'sh0be8f82c;
        7'b0110101 :  a = 32'sh0c3cf0a8;
        7'b0110110 :  a = 32'sh0c8dd9f8;
        7'b0110111 :  a = 32'sh0cdb9fe3;
        7'b0111000 :  a = 32'sh0d262ef6;
        7'b0111001 :  a = 32'sh0d6d7490;
        7'b0111010 :  a = 32'sh0db15ede;
        7'b0111011 :  a = 32'sh0df1dce6;
        7'b0111100 :  a = 32'sh0e2ede8a;
        7'b0111101 :  a = 32'sh0e685489;
        7'b0111110 :  a = 32'sh0e9e3087;
        7'b0111111 :  a = 32'sh0ed0650b;
        7'b1000000 :  a = 32'sh0efee58b;
        7'b1000001 :  a = 32'sh0f29a664;
        7'b1000010 :  a = 32'sh0f509ce9;
        7'b1000011 :  a = 32'sh0f73bf5a;
        7'b1000100 :  a = 32'sh0f9304f1;
        7'b1000101 :  a = 32'sh0fae65db;
        7'b1000110 :  a = 32'sh0fc5db40;
        7'b1000111 :  a = 32'sh0fd95f44;
        7'b1001000 :  a = 32'sh0fe8ed04;
        7'b1001001 :  a = 32'sh0ff4809f;
        7'b1001010 :  a = 32'sh0ffc172f;
        7'b1001011 :  a = 32'sh0fffaecf;
        7'b1001100 :  a = 32'sh0fff4698;
        7'b1001101 :  a = 32'sh0ffadea4;
        7'b1001110 :  a = 32'sh0ff2780f;
        7'b1001111 :  a = 32'sh0fe614f0;
        7'b1010000 :  a = 32'sh0fd5b862;
        7'b1010001 :  a = 32'sh0fc1667b;
        7'b1010010 :  a = 32'sh0fa9244f;
        7'b1010011 :  a = 32'sh0f8cf7ef;
        7'b1010100 :  a = 32'sh0f6ce865;
        7'b1010101 :  a = 32'sh0f48fdb6;
        7'b1010110 :  a = 32'sh0f2140dc;
        7'b1010111 :  a = 32'sh0ef5bbc6;
        7'b1011000 :  a = 32'sh0ec67955;
        7'b1011001 :  a = 32'sh0e938559;
        7'b1011010 :  a = 32'sh0e5cec90;
        7'b1011011 :  a = 32'sh0e22bc9e;
        7'b1011100 :  a = 32'sh0de50410;
        7'b1011101 :  a = 32'sh0da3d254;
        7'b1011110 :  a = 32'sh0d5f37b5;
        7'b1011111 :  a = 32'sh0d17455a;
        7'b1100000 :  a = 32'sh0ccc0d40;
        7'b1100001 :  a = 32'sh0c7da233;
        7'b1100010 :  a = 32'sh0c2c17ce;
        7'b1100011 :  a = 32'sh0bd78273;
        7'b1100100 :  a = 32'sh0b7ff748;
        7'b1100101 :  a = 32'sh0b258c2e;
        7'b1100110 :  a = 32'sh0ac857c0;
        7'b1100111 :  a = 32'sh0a68714a;
        7'b1101000 :  a = 32'sh0a05f0c6;
        7'b1101001 :  a = 32'sh09a0eed3;
        7'b1101010 :  a = 32'sh093984b1;
        7'b1101011 :  a = 32'sh08cfcc3a;
        7'b1101100 :  a = 32'sh0863dfdc;
        7'b1101101 :  a = 32'sh07f5da92;
        7'b1101110 :  a = 32'sh0785d7db;
        7'b1101111 :  a = 32'sh0713f3b8;
        7'b1110000 :  a = 32'sh06a04aa2;
        7'b1110001 :  a = 32'sh062af982;
        7'b1110010 :  a = 32'sh05b41dac;
        7'b1110011 :  a = 32'sh053bd4d6;
        7'b1110100 :  a = 32'sh04c23d11;
        7'b1110101 :  a = 32'sh044774c4;
        7'b1110110 :  a = 32'sh03cb9a9f;
        7'b1110111 :  a = 32'sh034ecd99;
        7'b1111000 :  a = 32'sh02d12ce4;
        7'b1111001 :  a = 32'sh0252d7e7;
        7'b1111010 :  a = 32'sh01d3ee38;
        7'b1111011 :  a = 32'sh01548f8f;
        7'b1111100 :  a = 32'sh00d4dbc4;
        7'b1111101 :  a = 32'sh0054f2c3;
        7'b1111110 :  a = 32'shffd4f487;
        7'b1111111 :  a = 32'shff55010c;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = 32'sh16a09e66;
        7'b0000001 :  b = 32'sh1752c7ca;
        7'b0000010 :  b = 32'sh17ff1c9b;
        7'b0000011 :  b = 32'sh18a571c5;
        7'b0000100 :  b = 32'sh19459db3;
        7'b0000101 :  b = 32'sh19df785b;
        7'b0000110 :  b = 32'sh1a72db48;
        7'b0000111 :  b = 32'sh1affa1a1;
        7'b0001000 :  b = 32'sh1b85a836;
        7'b0001001 :  b = 32'sh1c04cd86;
        7'b0001010 :  b = 32'sh1c7cf1c7;
        7'b0001011 :  b = 32'sh1cedf6f2;
        7'b0001100 :  b = 32'sh1d57c0c6;
        7'b0001101 :  b = 32'sh1dba34d1;
        7'b0001110 :  b = 32'sh1e153a76;
        7'b0001111 :  b = 32'sh1e68baf4;
        7'b0010000 :  b = 32'sh1eb4a16d;
        7'b0010001 :  b = 32'sh1ef8dae6;
        7'b0010010 :  b = 32'sh1f355652;
        7'b0010011 :  b = 32'sh1f6a0491;
        7'b0010100 :  b = 32'sh1f96d87a;
        7'b0010101 :  b = 32'sh1fbbc6d6;
        7'b0010110 :  b = 32'sh1fd8c66b;
        7'b0010111 :  b = 32'sh1fedcff9;
        7'b0011000 :  b = 32'sh1ffade3d;
        7'b0011001 :  b = 32'sh1fffedf5;
        7'b0011010 :  b = 32'sh1ffcfddc;
        7'b0011011 :  b = 32'sh1ff20eae;
        7'b0011100 :  b = 32'sh1fdf2326;
        7'b0011101 :  b = 32'sh1fc44001;
        7'b0011110 :  b = 32'sh1fa16bf6;
        7'b0011111 :  b = 32'sh1f76afba;
        7'b0100000 :  b = 32'sh1f4415fc;
        7'b0100001 :  b = 32'sh1f09ab62;
        7'b0100010 :  b = 32'sh1ec77e87;
        7'b0100011 :  b = 32'sh1e7d9ff5;
        7'b0100100 :  b = 32'sh1e2c2224;
        7'b0100101 :  b = 32'sh1dd31972;
        7'b0100110 :  b = 32'sh1d729c22;
        7'b0100111 :  b = 32'sh1d0ac253;
        7'b0101000 :  b = 32'sh1c9ba5f9;
        7'b0101001 :  b = 32'sh1c2562dc;
        7'b0101010 :  b = 32'sh1ba8168c;
        7'b0101011 :  b = 32'sh1b23e05b;
        7'b0101100 :  b = 32'sh1a98e156;
        7'b0101101 :  b = 32'sh1a073c3c;
        7'b0101110 :  b = 32'sh196f1576;
        7'b0101111 :  b = 32'sh18d0930c;
        7'b0110000 :  b = 32'sh182bdc9f;
        7'b0110001 :  b = 32'sh17811b5b;
        7'b0110010 :  b = 32'sh16d079ef;
        7'b0110011 :  b = 32'sh161a2484;
        7'b0110100 :  b = 32'sh155e48ac;
        7'b0110101 :  b = 32'sh149d155f;
        7'b0110110 :  b = 32'sh13d6bae8;
        7'b0110111 :  b = 32'sh130b6add;
        7'b0111000 :  b = 32'sh123b5811;
        7'b0111001 :  b = 32'sh1166b686;
        7'b0111010 :  b = 32'sh108dbb66;
        7'b0111011 :  b = 32'sh0fb09cec;
        7'b0111100 :  b = 32'sh0ecf9260;
        7'b0111101 :  b = 32'sh0dead404;
        7'b0111110 :  b = 32'sh0d029b05;
        7'b0111111 :  b = 32'sh0c172170;
        7'b1000000 :  b = 32'sh0b28a224;
        7'b1000001 :  b = 32'sh0a3758bd;
        7'b1000010 :  b = 32'sh0943818e;
        7'b1000011 :  b = 32'sh084d598b;
        7'b1000100 :  b = 32'sh07551e3d;
        7'b1000101 :  b = 32'sh065b0db1;
        7'b1000110 :  b = 32'sh055f666a;
        7'b1000111 :  b = 32'sh04626751;
        7'b1001000 :  b = 32'sh03644fa3;
        7'b1001001 :  b = 32'sh02655ee6;
        7'b1001010 :  b = 32'sh0165d4d5;
        7'b1001011 :  b = 32'sh0065f150;
        7'b1001100 :  b = 32'shff65f450;
        7'b1001101 :  b = 32'shfe661dd1;
        7'b1001110 :  b = 32'shfd66adca;
        7'b1001111 :  b = 32'shfc67e413;
        7'b1010000 :  b = 32'shfb6a005e;
        7'b1010001 :  b = 32'shfa6d4223;
        7'b1010010 :  b = 32'shf971e890;
        7'b1010011 :  b = 32'shf878327b;
        7'b1010100 :  b = 32'shf7805e4e;
        7'b1010101 :  b = 32'shf68aa9ff;
        7'b1010110 :  b = 32'shf59752f8;
        7'b1010111 :  b = 32'shf4a6960f;
        7'b1011000 :  b = 32'shf3b8af72;
        7'b1011001 :  b = 32'shf2cdda98;
        7'b1011010 :  b = 32'shf1e65236;
        7'b1011011 :  b = 32'shf102502c;
        7'b1011100 :  b = 32'shf0220d7b;
        7'b1011101 :  b = 32'shef45c231;
        7'b1011110 :  b = 32'shee6da560;
        7'b1011111 :  b = 32'shed99ed0e;
        7'b1100000 :  b = 32'sheccace28;
        7'b1100001 :  b = 32'shec007c76;
        7'b1100010 :  b = 32'sheb3b2a89;
        7'b1100011 :  b = 32'shea7b09b7;
        7'b1100100 :  b = 32'she9c04a05;
        7'b1100101 :  b = 32'she90b1a23;
        7'b1100110 :  b = 32'she85ba75c;
        7'b1100111 :  b = 32'she7b21d8b;
        7'b1101000 :  b = 32'she70ea713;
        7'b1101001 :  b = 32'she6716cd0;
        7'b1101010 :  b = 32'she5da960f;
        7'b1101011 :  b = 32'she54a4886;
        7'b1101100 :  b = 32'she4c0a847;
        7'b1101101 :  b = 32'she43dd7ba;
        7'b1101110 :  b = 32'she3c1f792;
        7'b1101111 :  b = 32'she34d26c6;
        7'b1110000 :  b = 32'she2df828b;
        7'b1110001 :  b = 32'she2792648;
        7'b1110010 :  b = 32'she21a2b94;
        7'b1110011 :  b = 32'she1c2aa2d;
        7'b1110100 :  b = 32'she172b7f3;
        7'b1110101 :  b = 32'she12a68e3;
        7'b1110110 :  b = 32'she0e9cf0f;
        7'b1110111 :  b = 32'she0b0fa9f;
        7'b1111000 :  b = 32'she07ff9c5;
        7'b1111001 :  b = 32'she056d8c4;
        7'b1111010 :  b = 32'she035a1e2;
        7'b1111011 :  b = 32'she01c5d6d;
        7'b1111100 :  b = 32'she00b11b6;
        7'b1111101 :  b = 32'she001c310;
        7'b1111110 :  b = 32'she00073cf;
        7'b1111111 :  b = 32'she0072446;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = 32'sh16a09e66;
        7'b0000001 :  c = 32'sh15e8ccf9;
        7'b0000010 :  c = 32'sh152b8176;
        7'b0000011 :  c = 32'sh1468eb2f;
        7'b0000100 :  c = 32'sh13a13ac8;
        7'b0000101 :  c = 32'sh12d4a22d;
        7'b0000110 :  c = 32'sh12035482;
        7'b0000111 :  c = 32'sh112d861a;
        7'b0001000 :  c = 32'sh10536c67;
        7'b0001001 :  c = 32'sh0f753def;
        7'b0001010 :  c = 32'sh0e93323c;
        7'b0001011 :  c = 32'sh0dad81d1;
        7'b0001100 :  c = 32'sh0cc46616;
        7'b0001101 :  c = 32'sh0bd81954;
        7'b0001110 :  c = 32'sh0ae8d69b;
        7'b0001111 :  c = 32'sh09f6d9ba;
        7'b0010000 :  c = 32'sh09025f31;
        7'b0010001 :  c = 32'sh080ba41c;
        7'b0010010 :  c = 32'sh0712e628;
        7'b0010011 :  c = 32'sh06186384;
        7'b0010100 :  c = 32'sh051c5ad0;
        7'b0010101 :  c = 32'sh041f0b0c;
        7'b0010110 :  c = 32'sh0320b38a;
        7'b0010111 :  c = 32'sh022193e0;
        7'b0011000 :  c = 32'sh0121ebd4;
        7'b0011001 :  c = 32'sh0021fb4e;
        7'b0011010 :  c = 32'shff220249;
        7'b0011011 :  c = 32'shfe2240c3;
        7'b0011100 :  c = 32'shfd22f6aa;
        7'b0011101 :  c = 32'shfc2463d0;
        7'b0011110 :  c = 32'shfb26c7d8;
        7'b0011111 :  c = 32'shfa2a6227;
        7'b0100000 :  c = 32'shf92f71d5;
        7'b0100001 :  c = 32'shf836359f;
        7'b0100010 :  c = 32'shf73eebd0;
        7'b0100011 :  c = 32'shf649d23b;
        7'b0100100 :  c = 32'shf5572624;
        7'b0100101 :  c = 32'shf4672436;
        7'b0100110 :  c = 32'shf37a086f;
        7'b0100111 :  c = 32'shf2900e15;
        7'b0101000 :  c = 32'shf1a96fa6;
        7'b0101001 :  c = 32'shf0c666c8;
        7'b0101010 :  c = 32'shefe72c3c;
        7'b0101011 :  c = 32'shef0bf7cf;
        7'b0101100 :  c = 32'shee35004e;
        7'b0101101 :  c = 32'shed627b75;
        7'b0101110 :  c = 32'shec949de4;
        7'b0101111 :  c = 32'shebcb9b12;
        7'b0110000 :  c = 32'sheb07a53e;
        7'b0110001 :  c = 32'shea48ed65;
        7'b0110010 :  c = 32'she98fa333;
        7'b0110011 :  c = 32'she8dbf4fb;
        7'b0110100 :  c = 32'she82e0fa7;
        7'b0110101 :  c = 32'she7861eaf;
        7'b0110110 :  c = 32'she6e44c0f;
        7'b0110111 :  c = 32'she648c03a;
        7'b0111000 :  c = 32'she5b3a213;
        7'b0111001 :  c = 32'she52516e1;
        7'b0111010 :  c = 32'she49d4245;
        7'b0111011 :  c = 32'she41c4633;
        7'b0111100 :  c = 32'she3a242ec;
        7'b0111101 :  c = 32'she32f56ed;
        7'b0111110 :  c = 32'she2c39ef2;
        7'b0111111 :  c = 32'she25f35e9;
        7'b1000000 :  c = 32'she20234eb;
        7'b1000001 :  c = 32'she1acb337;
        7'b1000010 :  c = 32'she15ec62e;
        7'b1000011 :  c = 32'she118814b;
        7'b1000100 :  c = 32'she0d9f61e;
        7'b1000101 :  c = 32'she0a3344b;
        7'b1000110 :  c = 32'she0744980;
        7'b1000111 :  c = 32'she04d4179;
        7'b1001000 :  c = 32'she02e25f7;
        7'b1001001 :  c = 32'she016fec2;
        7'b1001010 :  c = 32'she007d1a2;
        7'b1001011 :  c = 32'she000a263;
        7'b1001100 :  c = 32'she00172d1;
        7'b1001101 :  c = 32'she00a42b7;
        7'b1001110 :  c = 32'she01b0fe2;
        7'b1001111 :  c = 32'she033d61f;
        7'b1010000 :  c = 32'she0548f3c;
        7'b1010001 :  c = 32'she07d330b;
        7'b1010010 :  c = 32'she0adb762;
        7'b1010011 :  c = 32'she0e61023;
        7'b1010100 :  c = 32'she1262f36;
        7'b1010101 :  c = 32'she16e0494;
        7'b1010110 :  c = 32'she1bd7e48;
        7'b1010111 :  c = 32'she2148874;
        7'b1011000 :  c = 32'she2730d56;
        7'b1011001 :  c = 32'she2d8f54d;
        7'b1011010 :  c = 32'she34626e0;
        7'b1011011 :  c = 32'she3ba86c3;
        7'b1011100 :  c = 32'she435f7df;
        7'b1011101 :  c = 32'she4b85b58;
        7'b1011110 :  c = 32'she5419095;
        7'b1011111 :  c = 32'she5d1754b;
        7'b1100000 :  c = 32'she667e581;
        7'b1100001 :  c = 32'she704bb9b;
        7'b1100010 :  c = 32'she7a7d065;
        7'b1100011 :  c = 32'she850fb1a;
        7'b1100100 :  c = 32'she9001171;
        7'b1100101 :  c = 32'she9b4e7a4;
        7'b1100110 :  c = 32'shea6f5081;
        7'b1100111 :  c = 32'sheb2f1d6c;
        7'b1101000 :  c = 32'shebf41e74;
        7'b1101001 :  c = 32'shecbe225a;
        7'b1101010 :  c = 32'shed8cf69e;
        7'b1101011 :  c = 32'shee60678b;
        7'b1101100 :  c = 32'shef384047;
        7'b1101101 :  c = 32'shf0144add;
        7'b1101110 :  c = 32'shf0f4504a;
        7'b1101111 :  c = 32'shf1d81890;
        7'b1110000 :  c = 32'shf2bf6abc;
        7'b1110001 :  c = 32'shf3aa0cfc;
        7'b1110010 :  c = 32'shf497c4a9;
        7'b1110011 :  c = 32'shf5885655;
        7'b1110100 :  c = 32'shf67b85dd;
        7'b1110101 :  c = 32'shf7711678;
        7'b1110110 :  c = 32'shf868cac1;
        7'b1110111 :  c = 32'shf96264ce;
        7'b1111000 :  c = 32'shfa5da638;
        7'b1111001 :  c = 32'shfb5a5031;
        7'b1111010 :  c = 32'shfc582391;
        7'b1111011 :  c = 32'shfd56e0e2;
        7'b1111100 :  c = 32'shfe564878;
        7'b1111101 :  c = 32'shff561a79;
        7'b1111110 :  c = 32'sh005616f3;
        7'b1111111 :  c = 32'sh0155fde7;
        default    :  c = 'x;
    endcase

endmodule
